* C:\SPB_Data\eSim-Workspace\XOR\XOR.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 3/16/2021 10:29:54 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U1-Pad1_ Net-_U1-Pad3_ Net-_U3-Pad3_ nand_gate		
U2  Net-_U1-Pad3_ Net-_U1-Pad2_ Net-_U2-Pad3_ nand_gate		
U4  Net-_U3-Pad3_ Net-_U2-Pad3_ IN nand_gate		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ nand_gate		
v1  IN Net-_U1-Pad1_ pulse		
v2  Net-_U1-Pad2_ IN pulse		

.end
